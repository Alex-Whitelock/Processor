`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Rogue Squadron 
// Engineer: Alex, Logan,
// 
// Create Date:    12:51:14 10/24/2015 
// Design Name: 
// Module Name:    physical_tester 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module physical_tester(
    input clock,
    input reset,
    output [15:0] instruction
    );

//Test case was lost and will need to be re-written but we know that it is functioning due to test that were 
//written FPGA_REG_ALU_Display

endmodule
